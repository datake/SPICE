* kadai3-2-n16.cirs
***********************************************************************
* Set supply and library
***********************************************************************
.INCLUDE mos_model3
.options temp=27                * Nominal temperature
* Save results of simulation for viewing
.options post
***********************************************************************
* Define power supply
***********************************************************************
Vdd     Vdd     0       2.5
***********************************************************************
* Define Subcircuits
***********************************************************************
.subckt inv1 In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=32u
m2      Out In Vdd Vdd  cmosp l=0.25u w=64u
.ends

.subckt inv2 In Out Vdd
m1      Out In 0 0      cmosn l=0.25u w=4u
m2      Out In Vdd Vdd  cmosp l=0.25u w=2u
.ends


.subckt pi-model-wiring In Out 
R1	In	V1	20f
R2	V1	V2	40f
R3	V2	V3	40f
R4	V3	V4	40f
R5	V4	V5	40f
R6	V5	V6	40f
R7	V6	V7	40f
R8	V7	V8	40f
R9	V8	V9	40f
R10	V9	V10	40f
R11	V10	V11	40f
R12	V11	V12	40f
R13	V12	V13	40f
R14	V13	V14	40f
R15	V14	V15	40f
R16	V15	V16	20f




C1	V1	0	100p	
C2	V2	0   100p

.ends




***********************************************************************
* Stimulus
***********************************************************************
* Format of pulse input:
* pulse v_initial v_final t_delay t_rise t_fall t_pulsewidth t_period
V1     XA      0       PULSE(0 2.5 1ns 0.1ns 0.1ns 4ns 100ns)
V2      XB      0       PULSE(0 2.5 11ns 0.1ns 0.1ns 4ns 100ns)
V3      XC      0       PULSE(0 2.5 21ns 0.1ns 0.1ns 4ns 100ns)
V4      XD      0       PULSE(0 2.5 31ns 0.1ns 0.1ns 4ns 100ns)
***********************************************************************
* Top level simulation netlist
***********************************************************************
* ??? Add more of the netlist here
x1  XA  A Vdd inv
x2  XB  B Vdd inv
x3  XC  C Vdd inv
x4  XD  D Vdd inv

X1Nand   A B X1Nand_out Vdd NAND2
X2Nand   C D  X2Nand_out Vdd NAND2
 
X1Nor X1Nand_out X2Nand_out f Vdd NOR2



*xnand  A B C D NOUT Vdd NAND
*x5 NOUT F Vdd inv2
.tran .001ns 40ns
.plot TRAN V(A) V(B) V(C) V(D) V(vdd) V(XA) V(XB) V(XC) V(XD) V(NOUT) V(F)  V(x1nand_out)  V(x2nand_out)
***********************************************************************
* End of Deck
***********************************************************************
.end