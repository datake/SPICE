* kadai3-1-V1.cir
***********************************************************************
* Set supply and library
***********************************************************************
.INCLUDE mos_model3
.options temp=27                * Nominal temperature
* Save results of simulation for viewing
.options post
***********************************************************************
* Define power supply
***********************************************************************
Vdd     V0     0       PWL(On 0 0.1n 1)
***********************************************************************
* Top level simulation netlist
***********************************************************************
* ??? Add more of the netlist here
R1	V0	V1	100
C1	V1	0  300p
*x5 NOUT F Vdd inv2
.tran .001ns 300ns
.plot TRAN V(V1)
***********************************************************************
* End of Deck
***********************************************************************
.end